module clock_generator(
    clk,    //clock from crystal
    rst_n,  //active low reset
    clk_1,  //generated 1Hz clock
    clk_01,
    clk_100, //generated 100Hz clock
    clk_ctl //scan control
);
output clk_1;
output clk_01;
output clk_100;
output [1:0] clk_ctl;
input clk;
input rst_n;
reg clk_1;
reg clk_100;
reg clk_01;
reg [1:0] clk_ctl;

reg [26:0] count_50M, count_50M_next;
reg [26:0] count_5M, count_5M_next;
reg [26:0] count_500k, count_500k_next;
reg [26:0] count_100k, count_100k_next;

reg clk_1_next;
reg clk_100_next;
reg clk_01_next;
reg [1:0] clk_ctl_next;

//generate clock_ctl
always @*
    if (count_100k == 27'd100000)   //for display
    begin
        count_100k_next = 27'd0;
        clk_ctl_next = clk_ctl + 2'b1;
    end
    else
    begin
        count_100k_next = count_100k + 1'b1;
        clk_ctl_next = clk_ctl;
    end

always @(posedge clk or negedge rst_n)
    if (~rst_n)
    begin
        count_100k <= 27'd0;
        clk_ctl <= 2'b0;
    end
    else
    begin
        count_100k <= count_100k_next;
        clk_ctl <= clk_ctl_next;
    end

//generator clk_1 
always @*
    if (count_50M == 27'd50000000)
    begin
        count_50M_next = 27'd0;
        clk_1_next = ~clk_1;
    end
    else
    begin
        count_50M_next = count_50M + 1'b1;
        clk_1_next = clk_1;
    end

always @(posedge clk or negedge rst_n)
    if (~rst_n)
    begin
        count_50M <= 27'd0;
        clk_1 <= 1'b0;
    end
    else
    begin
        count_50M <= count_50M_next;
        clk_1 <= clk_1_next;
    end

//generator clk_01
always @*
    if (count_5M == 27'd5000000)
    begin
        count_5M_next = 27'd0;
        clk_01_next = ~clk_01;
    end
    else
    begin
        count_5M_next = count_5M + 1'b1;
        clk_01_next = clk_01;
    end

always @(posedge clk or negedge rst_n)
    if (~rst_n)
    begin
        count_5M <= 27'd0;
        clk_01 <= 1'b0;
    end
    else
    begin
        count_5M <= count_5M_next;
        clk_01 <= clk_01_next;
    end

//generator clk_100
always @*
    if (count_500k == 27'd500000)
    begin
        count_500k_next = 27'd0;
        clk_100_next = ~clk_100;
    end
    else
    begin
        count_500k_next = count_500k + 1'b1;
        clk_100_next = clk_100;
    end

always @(posedge clk or negedge rst_n)
    if (~rst_n)
    begin
        count_500k <= 27'd0;
        clk_100 <= 1'b0;
    end
    else
    begin
        count_500k <= count_500k_next;
        clk_100 <= clk_100_next;
    end
    
endmodule