module buzzer_control(
    clk,
    rst_n,
    vol,
    vol_minus,
    note_div_left,
    note_div_right,
    audio_left,
    audio_right
);
input clk;
input rst_n;
input [21:0] note_div_left, note_div_right;
input [15:0] vol, vol_minus;
output [15:0] audio_left;
output [15:0] audio_right;
reg [21:0] clk_cnt_next, clk_cnt;
reg [21:0] clk_cnt_2_next, clk_cnt_2;
reg b_clk, b_clk_next;
reg b_clk_2, b_clk_2_next;

always @(posedge clk or negedge rst_n)
    if (~rst_n)
    begin
        clk_cnt <= 22'd0;
        clk_cnt_2 <= 22'd0;
        b_clk <= 1'b0;
        b_clk_2 <= 1'b0;
    end
    else
    begin
        clk_cnt <= clk_cnt_next;
        clk_cnt_2 <= clk_cnt_2_next;
        b_clk <= b_clk_next;
        b_clk_2 <= b_clk_2_next;
    end

always @*
    if (clk_cnt == note_div_left)
    begin
        clk_cnt_next = 22'd0;
        b_clk_next = ~b_clk;
    end
    else
    begin
        clk_cnt_next = clk_cnt + 1'b1;
        b_clk_next = b_clk;
    end

always @*
    if (clk_cnt_2 == note_div_right)
    begin
        clk_cnt_2_next = 22'd0;
        b_clk_2_next = ~b_clk_2;
    end
    else
    begin
        clk_cnt_2_next = clk_cnt_2 + 1'b1;
        b_clk_2_next = b_clk_2;
    end

assign audio_left = (b_clk == 1'b0) ? vol_minus : vol;  //change the volume
assign audio_right = (b_clk_2 == 1'b0) ? vol_minus : vol; //change the volume

endmodule